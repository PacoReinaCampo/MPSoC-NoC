`include "peripheral_sequence_item.sv"
`include "peripheral_sequence.sv"
`include "peripheral_sequencer.sv"
`include "peripheral_driver.sv"
`include "peripheral_monitor.sv"
`include "peripheral_scoreboard.sv"
`include "peripheral_agent.sv"
`include "peripheral_enviroment.sv"